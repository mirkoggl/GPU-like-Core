fp_abs_inst : fp_abs PORT MAP (
		data	 => data_sig,
		result	 => result_sig
	);
